library verilog;
use verilog.vl_types.all;
entity SixteenBitAlu_vlg_vec_tst is
end SixteenBitAlu_vlg_vec_tst;
