library verilog;
use verilog.vl_types.all;
entity prob1_vlg_vec_tst is
end prob1_vlg_vec_tst;
