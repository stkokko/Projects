library verilog;
use verilog.vl_types.all;
entity OneBitAlu_vlg_vec_tst is
end OneBitAlu_vlg_vec_tst;
