library verilog;
use verilog.vl_types.all;
entity prob1_vlg_check_tst is
    port(
        h               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end prob1_vlg_check_tst;
